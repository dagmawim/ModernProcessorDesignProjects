library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity OR2 is
	port(x,y:in std_logic;z:out std_logic);
end OR2;
-- AND Operation on Two inputs
architecture behav of OR2 is
begin 
	z <= x or y;
end behav;